class msdap_scoreboard extends uvm_component;
  `uvm_component_utils(msdap_scoreboard)

  function new(string name = "msdap_scoreboard", uvm_component parent = null);
    super.new(name, parent);
  endfunction
endclass
