/proj/cad/library/asap7/asap7sc7p5t_28/techlef_misc/asap7_tech_1x_201209.lef