// Add config object here if needed
