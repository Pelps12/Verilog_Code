.SUBCKT SRAM2RW16x8 VDD VSS CE1 CE2 WEB1 WEB2 OEB1 OEB2 CSB1 CSB2 
+ A1[3] A1[2] A1[1] A1[0] A2[3] A2[2] A2[1] A2[0] 
+ I1[7] I1[6] I1[5] I1[4] I1[3] I1[2] I1[1] I1[0] 
+ I2[7] I2[6] I2[5] I2[4] I2[3] I2[2] I2[1] I2[0] 
+ O1[7] O1[6] O1[5] O1[4] O1[3] O1[2] O1[1] O1[0] 
+ O2[7] O2[6] O2[5] O2[4] O2[3] O2[2] O2[1] O2[0]
.ENDS SRAM2RW16x8

.SUBCKT SRAM1RW128x12 VDD VSS CE WEB OEB CSB A[6] A[5] A[4] A[3] A[2] A[1] A[0] 
+ I[11] I[10] I[9] I[8] I[7] I[6] I[5] I[4] I[3] I[2] I[1] I[0]
+ O[11] O[10] O[9] O[8] O[7] O[6] O[5] O[4] O[3] O[2] O[1] O[0]
.ENDS SRAM1RW128x12

.SUBCKT SRAM1RW256x8 VDD VSS CE WEB OEB CSB 
+ A[7] A[6] A[5] A[4] A[3] A[2] A[1] A[0]
+ I[7] I[6] I[5] I[4] I[3] I[2] I[1] I[0] 
+ O[7] O[6] O[5] O[4] O[3] O[2] O[1] O[0]
.ENDS SRAM1RW256x8


