/proj/cad/library/asap7/asap7sc7p5t_27/LEF/asap7sc7p5t_27_L_1x_201211.lef